// ============================================================================
//  Module: alu_slice4_nondep
// ----------------------------------------------------------------------------
//  Description:
//    4-bit ALU slice without inter-slice dependencies, designed specifically
//    for high-frequency operation on low-cost FPGAs.
//
//    This module is intended to be instantiated multiple times (e.g., 8 slices
//    for a 32-bit ALU). It follows a strict pipeline discipline and avoids
//    synthesis patterns that typically degrade Fmax on LUT-based fabrics.
//
//  Architectural Model:
//    - Explicit decode stage before execution
//    - One-hot operation signals pipelined alongside operands
//    - No carry propagation, no feedback loops
//    - Purely local logic per slice
//
//  Pipeline Stages:
//    Stage D (Decode / Register):
//      - Operands (a_in, b_in) are registered
//      - One-hot operation signals are registered
//      - Input validity (v_in) is captured
//
//    Stage X (Execute):
//      - All operations computed in parallel
//      - Result selected via logical masking (no wide multiplexers)
//
//    Stage W (Writeback / Register):
//      - Result registered
//      - Output validity asserted
//
//  FPGA-Oriented Design Techniques:
//    - Clock-enable inferred via if(v_in) / if(v_pipe)
//    - No combinational enable gating
//    - No wide multiplexers in the critical path
//    - No shared logic across slices
//    - Localized fanout and predictable placement
//
//  Assumptions:
//    - Only one do_* signal is asserted per valid instruction
//    - All do_* signals are generated by a prior decode stage
//    - do_* signals are stable when v_in is asserted
//
//  Notes:
//    - Registers are intentionally NOT reset
//    - Invalid cycles preserve previous data but deassert validity
//    - Designed for throughput and timing closure, not minimum area
//
// ============================================================================

module alu_slice4_nondep (
    input         clk,
    input         v_in,     // Input validity (from decode stage)

    input  [3:0]  a_in,     // Operand A
    input  [3:0]  b_in,     // Operand B

    // One-hot operation controls (from decode stage)
    input         do_and,
    input         do_or,
    input         do_xor,
    input         do_not,
    input         do_pass,

    output [3:0]  result,   // Registered result
    output        v_out     // Output validity
);

    // ------------------------------------------------------------------------
    // Stage D: Decode / Input Register Stage
    // Registers operands and one-hot operation signals.
    // This stage creates a hard pipeline boundary and limits fanout.
    // ------------------------------------------------------------------------

    reg [3:0] a_r;
    reg [3:0] b_r;

    reg do_and_r;
    reg do_or_r;
    reg do_xor_r;
    reg do_not_r;
    reg do_pass_r;

    reg v_pipe;

    always @(posedge clk) begin
        if (v_in) begin
            a_r       <= a_in;
            b_r       <= b_in;

            do_and_r  <= do_and;
            do_or_r   <= do_or;
            do_xor_r  <= do_xor;
            do_not_r  <= do_not;
            do_pass_r <= do_pass;

            v_pipe    <= 1'b1;
        end else begin
            v_pipe    <= 1'b0;
        end
    end

    // ------------------------------------------------------------------------
    // Stage X: Execute (Combinational, fully parallel)
    // All operations are computed unconditionally.
    // Selection is done via logical masking (no multiplexers).
    // ------------------------------------------------------------------------

    wire [3:0] and_res  = a_r & b_r;
    wire [3:0] or_res   = a_r | b_r;
    wire [3:0] xor_res  = a_r ^ b_r;
    wire [3:0] not_res  = ~a_r;
    wire [3:0] pass_res = a_r;

    wire [3:0] result_c =
          ({4{do_and_r }} & and_res )
        | ({4{do_or_r  }} & or_res  )
        | ({4{do_xor_r }} & xor_res )
        | ({4{do_not_r }} & not_res )
        | ({4{do_pass_r}} & pass_res);

    // ------------------------------------------------------------------------
    // Stage W: Writeback / Output Register Stage
    // Registers the result and propagates validity.
    // ------------------------------------------------------------------------

    reg [3:0] result_r;
    reg       v_out_r;

    always @(posedge clk) begin
        if (v_pipe) begin
            result_r <= result_c;
            v_out_r  <= 1'b1;
        end else begin
            v_out_r  <= 1'b0;
        end
    end

    assign result = result_r;
    assign v_out  = v_out_r;

endmodule
